// Create a 100-bit binary adder. The adder adds two 100-bit numbers and a carry-in to produce a 100-bit sum and carry out.
module top_module( 
    input [99:0] a, b,
    input cin,
    output cout,
    output [99:0] sum );
	assign {cout, ss} = a + b + cin;
endmodule
